module inverter(in, out);

input in;
output wire out;

assign out = ~in; 

endmodule
